module fadd(a,b,out);
endmodule
