//assign kgp to each c
module kgp(a,b,c);
input a,b;
output [1:0]c;
wire [1:0]k,g,p;
reg [1:0]c;
assign k=2'b00;
assign p=2'b10;
assign g=2'b11;
always@(a or b)
begin
c=(a==b)?(a==1)?g:k:p;
end
endmodule



module padd(a,b,c);
input [63:0] a,b ;
output [129:0] c;
assign c[1:0]=2'b00; 
kgp t0(a[0],b[0],c[3:2]);
kgp t1(a[1],b[1],c[5:4]);
kgp t2(a[2],b[2],c[7:6]);
kgp t3(a[3],b[3],c[9:8]);
kgp t4(a[4],b[4],c[11:10]);
kgp t5(a[5],b[5],c[13:12]);
kgp t6(a[6],b[6],c[15:14]);
kgp t7(a[7],b[7],c[17:16]);
kgp t8(a[8],b[8],c[19:18]);
kgp t9(a[9],b[9],c[21:20]);
kgp t10(a[10],b[10],c[23:22]);
kgp t11(a[11],b[11],c[25:24]);
kgp t12(a[12],b[12],c[27:26]);
kgp t13(a[13],b[13],c[29:28]); 
kgp t14(a[14],b[14],c[31:30]); 
kgp t15(a[15],b[15],c[33:32]); 
kgp t16(a[16],b[16],c[35:34]);
kgp t17(a[17],b[17],c[37:36]);
kgp t18(a[18],b[18],c[39:38]);
kgp t19(a[19],b[19],c[41:40]);
kgp t20(a[20],b[20],c[43:42]);
kgp t21(a[21],b[21],c[45:44]);
kgp t22(a[22],b[22],c[47:46]);
kgp t23(a[23],b[23],c[49:48]);
kgp t24(a[24],b[24],c[51:50]);
kgp t25(a[25],b[25],c[53:52]);
kgp t26(a[26],b[26],c[55:54]);
kgp t27(a[27],b[27],c[57:56]);
kgp t28(a[28],b[28],c[59:58]);
kgp t29(a[29],b[29],c[61:60]); 
kgp t30(a[30],b[30],c[63:62]); 
kgp t31(a[31],b[31],c[65:64]); 
kgp t32(a[32],b[32],c[67:66]);
kgp t33(a[33],b[33],c[69:68]);
kgp t34(a[34],b[34],c[71:70]);
kgp t35(a[35],b[35],c[73:72]);
kgp t36(a[36],b[36],c[75:74]);
kgp t37(a[37],b[37],c[77:76]);
kgp t38(a[38],b[38],c[79:78]);
kgp t39(a[39],b[39],c[81:80]);
kgp t40(a[40],b[40],c[83:82]);
kgp t41(a[41],b[41],c[85:84]);
kgp t42(a[42],b[42],c[87:86]);
kgp t43(a[43],b[43],c[89:88]);
kgp t44(a[44],b[44],c[91:90]);
kgp t45(a[45],b[45],c[93:92]); 
kgp t46(a[46],b[46],c[95:94]); 
kgp t47(a[47],b[47],c[97:96]);
kgp t48(a[48],b[48],c[99:98]);
kgp t49(a[49],b[49],c[101:100]);
kgp t50(a[50],b[50],c[103:102]);
kgp t51(a[51],b[51],c[105:104]);
kgp t52(a[52],b[52],c[107:106]);
kgp t53(a[53],b[53],c[109:108]);
kgp t54(a[54],b[54],c[111:110]);
kgp t55(a[55],b[55],c[113:112]);
kgp t56(a[56],b[56],c[115:114]);
kgp t57(a[57],b[57],c[117:116]);
kgp t58(a[58],b[58],c[119:118]);
kgp t59(a[59],b[59],c[121:120]);
kgp t60(a[60],b[60],c[123:122]);
kgp t61(a[61],b[61],c[125:124]); 
kgp t62(a[62],b[62],c[127:126]); 
kgp t63(a[63],b[63],c[129:128]); 
endmodule 


module padd1(x,y);
input [129:0]x;
output [129:0]y;
reg [129:0]y;
reg [2:0]p;
always@(x)
begin
p=2'b10;
y=x;
y[129:128]=(x[129:128]==p)?x[127:126]:y[129:128];
y[127:126]=(x[127:126]==p)?x[125:124]:y[127:126];
y[125:124]=(x[125:124]==p)?x[123:122]:y[125:124];
y[123:122]=(x[123:122]==p)?x[121:120]:y[123:122];
y[121:120]=(x[121:120]==p)?x[119:118]:y[121:120];
y[119:118]=(x[119:118]==p)?x[117:116]:y[119:118];
y[117:116]=(x[117:116]==p)?x[115:114]:y[117:116];
y[115:114]=(x[115:114]==p)?x[113:112]:y[115:114];
y[113:112]=(x[113:112]==p)?x[111:110]:y[113:112];
y[111:110]=(x[111:110]==p)?x[109:108]:y[111:110];
y[109:108]=(x[109:108]==p)?x[107:106]:y[109:108];
y[107:106]=(x[107:106]==p)?x[105:104]:y[107:106];
y[105:104]=(x[105:104]==p)?x[103:102]:y[105:104];
y[103:102]=(x[103:102]==p)?x[101:100]:y[103:102];
y[101:100]=(x[101:100]==p)?x[99:98]:y[101:100];
y[99:98]=(x[99:98]==p)?x[97:96]:y[99:98];
y[97:96]=(x[97:96]==p)?x[95:94]:y[97:96];
y[95:94]=(x[95:94]==p)?x[93:92]:y[95:94];
y[93:92]=(x[93:92]==p)?x[91:90]:y[93:92];
y[91:90]=(x[91:90]==p)?x[89:88]:y[91:90];
y[89:88]=(x[89:88]==p)?x[87:86]:y[89:88];
y[87:86]=(x[87:86]==p)?x[85:84]:y[87:86];
y[85:84]=(x[85:84]==p)?x[83:82]:y[85:84];
y[83:82]=(x[83:82]==p)?x[81:80]:y[83:82];
y[81:80]=(x[81:80]==p)?x[79:78]:y[81:80];
y[79:78]=(x[79:78]==p)?x[77:76]:y[79:78];
y[77:76]=(x[77:76]==p)?x[75:74]:y[77:76];
y[75:74]=(x[75:74]==p)?x[73:72]:y[75:74];
y[73:72]=(x[73:72]==p)?x[71:70]:y[73:72];
y[71:70]=(x[71:70]==p)?x[69:68]:y[71:70];
y[69:68]=(x[69:68]==p)?x[67:66]:y[69:68];
y[67:66]=(x[67:66]==p)?x[65:64]:y[67:66];
y[65:64]=(x[65:64]==p)?x[63:62]:y[65:64];
y[63:22]=(x[63:62]==p)?x[61:60]:y[63:22];
y[61:60]=(x[61:60]==p)?x[59:58]:y[61:60];
y[59:58]=(x[59:58]==p)?x[57:56]:y[59:58];
y[57:56]=(x[57:56]==p)?x[55:54]:y[57:56];
y[55:54]=(x[55:54]==p)?x[53:52]:y[55:54];
y[53:52]=(x[53:52]==p)?x[51:50]:y[53:52];
y[51:50]=(x[51:50]==p)?x[49:48]:y[51:50];
y[49:48]=(x[49:48]==p)?x[47:46]:y[49:48];
y[47:46]=(x[47:46]==p)?x[45:44]:y[47:46];
y[45:44]=(x[45:44]==p)?x[43:42]:y[45:44];
y[43:42]=(x[43:42]==p)?x[41:40]:y[43:42];
y[41:40]=(x[41:40]==p)?x[39:38]:y[41:40];
y[39:38]=(x[39:38]==p)?x[37:36]:y[39:38];
y[37:36]=(x[37:36]==p)?x[35:34]:y[37:36];
y[35:34]=(x[35:34]==p)?x[33:32]:y[35:34];
y[33:32]=(x[33:32]==p)?x[31:30]:y[33:32];
y[31:30]=(x[31:30]==p)?x[29:28]:y[31:30];
y[29:28]=(x[29:28]==p)?x[27:26]:y[29:28];
y[27:26]=(x[27:26]==p)?x[25:24]:y[27:26];
y[25:24]=(x[25:24]==p)?x[23:22]:y[25:24];
y[23:22]=(x[23:22]==p)?x[21:20]:y[23:22];
y[21:20]=(x[21:20]==p)?x[19:18]:y[21:20];
y[19:18]=(x[19:18]==p)?x[17:16]:y[19:18];
y[17:16]=(x[17:16]==p)?x[15:14]:y[17:16];
y[15:14]=(x[15:14]==p)?x[13:12]:y[15:14];
y[13:12]=(x[13:12]==p)?x[11:10]:y[13:12];
y[11:10]=(x[11:10]==p)?x[9:8]:y[11:10];
y[9:8]=(x[9:8]==p)?x[7:6]:y[9:8];
y[7:6]=(x[7:6]==p)?x[5:4]:y[7:6];
y[5:4]=(x[5:4]==p)?x[3:2]:y[5:4];
y[3:2]=(x[3:2]==p)?x[1:0]:y[3:2];
end
endmodule

module padd2(x,y);
input [129:0]x;
output [129:0]y;
reg [129:0]y;
reg [2:0]p;
always@(x)
begin
p=2'b10;
y=x;
y[129:128]=(x[129:128]==p)?x[125:124]:y[129:128];
y[127:126]=(x[127:126]==p)?x[123:122]:y[127:126];
y[125:124]=(x[125:124]==p)?x[121:120]:y[125:124];
y[123:122]=(x[123:122]==p)?x[119:118]:y[123:122];
y[121:120]=(x[121:120]==p)?x[117:116]:y[121:120];
y[119:118]=(x[119:118]==p)?x[115:114]:y[119:118];
y[117:116]=(x[117:116]==p)?x[113:112]:y[117:116];
y[115:114]=(x[115:114]==p)?x[111:110]:y[115:114];
y[113:112]=(x[113:112]==p)?x[109:108]:y[113:112];
y[111:110]=(x[111:110]==p)?x[107:106]:y[111:110];
y[109:108]=(x[109:108]==p)?x[105:104]:y[109:108];
y[107:106]=(x[107:106]==p)?x[103:102]:y[107:106];
y[105:104]=(x[105:104]==p)?x[101:100]:y[105:104];
y[103:102]=(x[103:102]==p)?x[99:98]:y[103:102];
y[101:100]=(x[101:100]==p)?x[97:96]:y[101:100];
y[99:98]=(x[99:98]==p)?x[95:94]:y[99:98];
y[97:96]=(x[97:96]==p)?x[93:92]:y[97:97];
y[95:94]=(x[95:94]==p)?x[91:90]:y[95:94];
y[93:92]=(x[93:92]==p)?x[89:88]:y[93:92];
y[91:90]=(x[91:90]==p)?x[87:86]:y[91:90];
y[89:88]=(x[89:88]==p)?x[85:84]:y[89:88];
y[87:86]=(x[87:86]==p)?x[83:82]:y[87:86];
y[85:84]=(x[85:84]==p)?x[81:80]:y[85:84];
y[83:82]=(x[83:82]==p)?x[79:78]:y[83:82];
y[81:80]=(x[81:80]==p)?x[77:76]:y[81:80];
y[79:78]=(x[79:78]==p)?x[75:74]:y[79:78];
y[77:76]=(x[77:76]==p)?x[73:72]:y[77:76];
y[75:74]=(x[75:74]==p)?x[71:70]:y[75:74];
y[73:72]=(x[73:72]==p)?x[69:68]:y[73:72];
y[71:70]=(x[71:70]==p)?x[67:66]:y[71:70];
y[69:68]=(x[69:68]==p)?x[65:64]:y[69:68];
y[67:66]=(x[67:66]==p)?x[63:62]:y[67:66];
y[65:64]=(x[65:64]==p)?x[61:60]:y[65:64];
y[63:62]=(x[63:62]==p)?x[59:58]:y[63:62];
y[61:60]=(x[61:60]==p)?x[57:56]:y[61:60];
y[59:58]=(x[59:58]==p)?x[55:54]:y[59:58];
y[57:56]=(x[57:56]==p)?x[53:52]:y[57:56];
y[55:54]=(x[55:54]==p)?x[51:50]:y[55:54];
y[53:52]=(x[53:52]==p)?x[49:48]:y[53:52];
y[51:50]=(x[51:50]==p)?x[47:46]:y[51:50];
y[49:48]=(x[49:48]==p)?x[45:44]:y[49:48];
y[47:46]=(x[47:46]==p)?x[43:42]:y[47:46];
y[45:44]=(x[45:44]==p)?x[41:40]:y[45:44];
y[43:42]=(x[43:42]==p)?x[39:38]:y[43:42];
y[41:40]=(x[41:40]==p)?x[37:36]:y[41:40];
y[39:38]=(x[39:38]==p)?x[35:34]:y[39:38];
y[37:36]=(x[37:36]==p)?x[33:32]:y[37:36];
y[35:34]=(x[35:34]==p)?x[31:30]:y[35:34];
y[33:32]=(x[33:32]==p)?x[29:28]:y[33:32];
y[31:30]=(x[31:30]==p)?x[27:26]:y[31:30];
y[29:28]=(x[29:28]==p)?x[25:24]:y[29:28];
y[27:26]=(x[27:26]==p)?x[23:22]:y[27:26];
y[25:24]=(x[25:24]==p)?x[21:20]:y[25:24];
y[23:22]=(x[23:22]==p)?x[19:18]:y[23:22];
y[21:20]=(x[21:20]==p)?x[17:16]:y[21:20];
y[19:18]=(x[19:18]==p)?x[15:14]:y[19:18];
y[17:16]=(x[17:16]==p)?x[13:12]:y[17:16];
y[15:14]=(x[15:14]==p)?x[11:10]:y[15:14];
y[13:12]=(x[13:12]==p)?x[9:8]:y[13:12];
y[11:10]=(x[11:10]==p)?x[7:6]:y[11:10];
y[9:8]=(x[9:8]==p)?x[5:4]:y[9:8];
y[7:6]=(x[7:6]==p)?x[3:2]:y[7:6];
y[5:4]=(x[5:4]==p)?x[1:0]:y[5:4];
end
endmodule


module padd3(x,y);
input [129:0]x;
output [129:0]y;
reg [129:0]y;
reg [2:0]p;
always@(x)
begin
p=2'b10;
y=x;
y[129:128]=(x[129:128]==p)?x[121:120]:y[129:128];
y[127:126]=(x[127:126]==p)?x[119:118]:y[127:126];
y[125:124]=(x[125:124]==p)?x[117:116]:y[125:124];
y[123:122]=(x[123:122]==p)?x[115:114]:y[123:122];
y[121:120]=(x[121:120]==p)?x[113:112]:y[121:120];
y[119:118]=(x[119:118]==p)?x[111:110]:y[119:118];
y[117:116]=(x[117:116]==p)?x[109:108]:y[117:116];
y[115:114]=(x[115:114]==p)?x[107:106]:y[115:114];
y[113:112]=(x[113:112]==p)?x[105:104]:y[113:112];
y[111:110]=(x[111:110]==p)?x[103:102]:y[111:110];
y[109:108]=(x[109:108]==p)?x[101:100]:y[109:108];
y[107:106]=(x[107:106]==p)?x[99:98]:y[107:106];
y[105:104]=(x[105:104]==p)?x[97:96]:y[105:104];
y[103:102]=(x[103:102]==p)?x[95:94]:y[103:102];
y[101:100]=(x[101:100]==p)?x[93:92]:y[101:100];
y[99:98]=(x[99:98]==p)?x[91:90]:y[99:98];
y[97:97]=(x[97:96]==p)?x[89:88]:y[97:97];
y[95:94]=(x[95:94]==p)?x[87:86]:y[95:94];
y[93:92]=(x[93:92]==p)?x[85:84]:y[93:92];
y[91:90]=(x[91:90]==p)?x[83:82]:y[91:90];
y[89:88]=(x[89:88]==p)?x[81:80]:y[89:88];
y[87:86]=(x[87:86]==p)?x[79:78]:y[87:86];
y[85:84]=(x[85:84]==p)?x[77:76]:y[85:84];
y[83:82]=(x[83:82]==p)?x[75:74]:y[83:82];
y[81:80]=(x[81:80]==p)?x[73:72]:y[81:80];
y[79:78]=(x[79:78]==p)?x[71:70]:y[79:78];
y[77:76]=(x[77:76]==p)?x[69:68]:y[77:76];
y[75:74]=(x[75:74]==p)?x[67:66]:y[75:74];
y[73:72]=(x[73:72]==p)?x[65:64]:y[73:72];
y[71:70]=(x[71:70]==p)?x[63:62]:y[71:70];
y[69:68]=(x[69:68]==p)?x[61:60]:y[69:68];
y[67:66]=(x[67:66]==p)?x[59:58]:y[67:66];
y[65:64]=(x[65:64]==p)?x[57:56]:y[65:64];
y[63:62]=(x[63:62]==p)?x[55:54]:y[63:62];
y[61:60]=(x[61:60]==p)?x[53:52]:y[61:60];
y[59:58]=(x[59:58]==p)?x[51:50]:y[59:58];
y[57:56]=(x[57:56]==p)?x[49:48]:y[57:56];
y[55:54]=(x[55:54]==p)?x[47:46]:y[55:54];
y[53:52]=(x[53:52]==p)?x[45:44]:y[53:52];
y[51:50]=(x[51:50]==p)?x[43:42]:y[51:50];
y[49:48]=(x[49:48]==p)?x[41:40]:y[49:48];
y[47:46]=(x[47:46]==p)?x[39:38]:y[47:46];
y[45:44]=(x[45:44]==p)?x[37:36]:y[45:44];
y[43:42]=(x[43:42]==p)?x[35:34]:y[43:42];
y[41:40]=(x[41:40]==p)?x[33:32]:y[41:40];
y[39:38]=(x[39:38]==p)?x[31:30]:y[39:38];
y[37:36]=(x[37:36]==p)?x[29:28]:y[37:36];
y[35:34]=(x[35:34]==p)?x[27:26]:y[35:34];
y[33:32]=(x[33:32]==p)?x[25:24]:y[33:32];
y[31:30]=(x[31:30]==p)?x[23:22]:y[31:30];
y[29:28]=(x[29:28]==p)?x[21:20]:y[29:28];
y[27:26]=(x[27:26]==p)?x[19:18]:y[27:26];
y[25:24]=(x[25:24]==p)?x[17:16]:y[25:24];
y[23:22]=(x[23:22]==p)?x[15:14]:y[23:22];
y[21:20]=(x[21:20]==p)?x[13:12]:y[21:20];
y[19:18]=(x[19:18]==p)?x[11:10]:y[19:18];
y[17:16]=(x[17:16]==p)?x[9:8]:y[17:16];
y[15:14]=(x[15:14]==p)?x[7:6]:y[15:14];
y[13:12]=(x[13:12]==p)?x[5:4]:y[13:12];
y[11:10]=(x[11:10]==p)?x[3:2]:y[11:10];
y[9:8]=(x[9:8]==p)?x[1:0]:y[9:8];
end
endmodule

module padd4(x,y);
input [129:0]x;
output [129:0]y;
reg [129:0]y;
reg [2:0]p;
always@(x)
begin
p=2'b10;
y=x;
y[129:128]=(x[129:128]==p)?x[113:112]:y[129:128];
y[127:126]=(x[127:126]==p)?x[111:110]:y[127:126];
y[125:124]=(x[125:124]==p)?x[109:108]:y[125:124];
y[123:122]=(x[123:122]==p)?x[107:106]:y[123:122];
y[121:120]=(x[121:120]==p)?x[105:104]:y[121:120];
y[119:118]=(x[119:118]==p)?x[103:102]:y[119:118];
y[117:116]=(x[117:116]==p)?x[101:100]:y[117:116];
y[115:114]=(x[115:114]==p)?x[99:98]:y[115:114];
y[113:112]=(x[113:112]==p)?x[97:96]:y[113:112];
y[111:110]=(x[111:110]==p)?x[95:94]:y[111:110];
y[109:108]=(x[109:108]==p)?x[93:92]:y[109:108];
y[107:106]=(x[107:106]==p)?x[91:90]:y[107:106];
y[105:104]=(x[105:104]==p)?x[89:88]:y[105:104];
y[103:102]=(x[103:102]==p)?x[87:86]:y[103:102];
y[101:100]=(x[101:100]==p)?x[85:84]:y[101:100];
y[99:98]=(x[99:98]==p)?x[83:82]:y[99:98];
y[97:97]=(x[97:96]==p)?x[81:80]:y[97:97];
y[95:94]=(x[95:94]==p)?x[79:78]:y[95:94];
y[93:92]=(x[93:92]==p)?x[77:76]:y[93:92];
y[91:90]=(x[91:90]==p)?x[75:74]:y[91:90];
y[89:88]=(x[89:88]==p)?x[73:72]:y[89:88];
y[87:86]=(x[87:86]==p)?x[71:70]:y[87:86];
y[85:84]=(x[85:84]==p)?x[69:68]:y[85:84];
y[83:82]=(x[83:82]==p)?x[67:66]:y[83:82];
y[81:80]=(x[81:80]==p)?x[65:64]:y[81:80];
y[79:78]=(x[79:78]==p)?x[63:62]:y[79:78];
y[77:76]=(x[77:76]==p)?x[61:60]:y[77:76];
y[75:74]=(x[75:74]==p)?x[59:58]:y[75:74];
y[73:72]=(x[73:72]==p)?x[57:56]:y[73:72];
y[71:70]=(x[71:70]==p)?x[55:54]:y[71:70];
y[69:68]=(x[69:68]==p)?x[53:52]:y[69:68];
y[67:66]=(x[67:66]==p)?x[51:50]:y[67:66];
y[65:64]=(x[65:64]==p)?x[49:48]:y[65:64];
y[63:62]=(x[63:62]==p)?x[47:46]:y[63:62];
y[61:60]=(x[61:60]==p)?x[45:44]:y[61:60];
y[59:58]=(x[59:58]==p)?x[43:42]:y[59:58];
y[57:56]=(x[57:56]==p)?x[41:40]:y[57:56];
y[55:54]=(x[55:54]==p)?x[39:38]:y[55:54];
y[53:52]=(x[53:52]==p)?x[37:36]:y[53:52];
y[51:50]=(x[51:50]==p)?x[35:34]:y[51:50];
y[49:48]=(x[49:48]==p)?x[33:32]:y[49:48];
y[47:46]=(x[47:46]==p)?x[31:30]:y[47:46];
y[45:44]=(x[45:44]==p)?x[29:28]:y[45:44];
y[43:42]=(x[43:42]==p)?x[27:26]:y[43:42];
y[41:40]=(x[41:40]==p)?x[25:24]:y[41:40];
y[39:38]=(x[39:38]==p)?x[23:22]:y[39:38];
y[37:36]=(x[37:36]==p)?x[21:20]:y[37:36];
y[35:34]=(x[35:34]==p)?x[19:18]:y[35:34];
y[33:32]=(x[33:32]==p)?x[17:16]:y[33:32];
y[31:30]=(x[31:30]==p)?x[15:14]:y[31:30];
y[29:28]=(x[29:28]==p)?x[13:12]:y[29:28];
y[27:26]=(x[27:26]==p)?x[11:10]:y[27:26];
y[25:24]=(x[25:24]==p)?x[9:8]:y[25:24];
y[23:22]=(x[23:22]==p)?x[7:6]:y[23:22];
y[21:20]=(x[21:20]==p)?x[5:4]:y[21:20];
y[19:18]=(x[19:18]==p)?x[3:2]:y[19:18];
y[17:16]=(x[17:16]==p)?x[1:0]:y[17:16];
end
endmodule


module padd5(x,y);
input [129:0]x;
output [129:0]y;
reg [129:0]y;
reg [2:0]p;
always@(x)
begin
p=2'b10;
y=x;
y[129:128]=(x[129:128]==p)?x[97:96]:y[129:128];
y[127:126]=(x[127:126]==p)?x[95:94]:y[127:126];
y[125:124]=(x[125:124]==p)?x[93:92]:y[125:124];
y[123:122]=(x[123:122]==p)?x[91:90]:y[123:122];
y[121:120]=(x[121:120]==p)?x[89:88]:y[121:120];
y[119:118]=(x[119:118]==p)?x[87:86]:y[119:118];
y[117:116]=(x[117:116]==p)?x[85:84]:y[117:116];
y[115:114]=(x[115:114]==p)?x[83:82]:y[115:114];
y[113:112]=(x[113:112]==p)?x[81:80]:y[113:112];
y[111:110]=(x[111:110]==p)?x[79:78]:y[111:110];
y[109:108]=(x[109:108]==p)?x[77:76]:y[109:108];
y[107:106]=(x[107:106]==p)?x[75:74]:y[107:106];
y[105:104]=(x[105:104]==p)?x[73:72]:y[105:104];
y[103:102]=(x[103:102]==p)?x[71:70]:y[103:102];
y[101:100]=(x[101:100]==p)?x[69:68]:y[101:100];
y[99:98]=(x[99:98]==p)?x[67:66]:y[99:98];
y[97:97]=(x[97:96]==p)?x[65:64]:y[97:97];
y[95:94]=(x[95:94]==p)?x[63:62]:y[95:94];
y[93:92]=(x[93:92]==p)?x[61:60]:y[93:92];
y[91:90]=(x[91:90]==p)?x[59:58]:y[91:90];
y[89:88]=(x[89:88]==p)?x[57:56]:y[89:88];
y[87:86]=(x[87:86]==p)?x[55:54]:y[87:86];
y[85:84]=(x[85:84]==p)?x[53:52]:y[85:84];
y[83:82]=(x[83:82]==p)?x[51:50]:y[83:82];
y[81:80]=(x[81:80]==p)?x[49:48]:y[81:80];
y[79:78]=(x[79:78]==p)?x[47:46]:y[79:78];
y[77:76]=(x[77:76]==p)?x[45:44]:y[77:76];
y[75:74]=(x[75:74]==p)?x[43:42]:y[75:74];
y[73:72]=(x[73:72]==p)?x[41:40]:y[73:72];
y[71:70]=(x[71:70]==p)?x[39:38]:y[71:70];
y[69:68]=(x[69:68]==p)?x[37:36]:y[69:68];
y[67:66]=(x[67:66]==p)?x[35:34]:y[67:66];
y[65:64]=(x[65:64]==p)?x[33:32]:y[65:64];
y[63:22]=(x[63:62]==p)?x[31:30]:y[63:22];
y[61:60]=(x[61:60]==p)?x[29:28]:y[61:60];
y[59:58]=(x[59:58]==p)?x[27:26]:y[59:58];
y[57:56]=(x[57:56]==p)?x[25:24]:y[57:56];
y[55:54]=(x[55:54]==p)?x[23:22]:y[55:54];
y[53:52]=(x[53:52]==p)?x[21:20]:y[53:52];
y[51:50]=(x[51:50]==p)?x[19:18]:y[51:50];
y[49:48]=(x[49:48]==p)?x[17:16]:y[49:48];
y[47:46]=(x[47:46]==p)?x[15:14]:y[47:46];
y[45:44]=(x[45:44]==p)?x[13:12]:y[45:44];
y[43:42]=(x[43:42]==p)?x[11:10]:y[43:42];
y[41:40]=(x[41:40]==p)?x[9:8]:y[41:40];
y[39:38]=(x[39:38]==p)?x[7:6]:y[39:38];
y[37:36]=(x[37:36]==p)?x[5:4]:y[37:36];
y[35:34]=(x[35:34]==p)?x[3:2]:y[35:34];
y[33:32]=(x[33:32]==p)?x[1:0]:y[33:32];
end
endmodule



module padd6(x,y);
input [129:0]x;
output [129:0]y;
reg [129:0]y;
reg [2:0]p;
always@(x)
begin
p=2'b10;
y=x;
y[129:128]=(x[129:128]==p)?x[65:64]:y[129:128];
y[127:126]=(x[127:126]==p)?x[63:62]:y[127:126];
y[125:124]=(x[125:124]==p)?x[61:60]:y[125:124];
y[123:122]=(x[123:122]==p)?x[59:58]:y[123:122];
y[121:120]=(x[121:120]==p)?x[57:56]:y[121:120];
y[119:118]=(x[119:118]==p)?x[55:54]:y[119:118];
y[117:116]=(x[117:116]==p)?x[53:52]:y[117:116];
y[115:114]=(x[115:114]==p)?x[51:50]:y[115:114];
y[113:112]=(x[113:112]==p)?x[49:48]:y[113:112];
y[111:110]=(x[111:110]==p)?x[47:46]:y[111:110];
y[109:108]=(x[109:108]==p)?x[45:44]:y[109:108];
y[107:106]=(x[107:106]==p)?x[43:42]:y[107:106];
y[105:104]=(x[105:104]==p)?x[41:40]:y[105:104];
y[103:102]=(x[103:102]==p)?x[39:38]:y[103:102];
y[101:100]=(x[101:100]==p)?x[37:36]:y[101:100];
y[99:98]=(x[99:98]==p)?x[35:34]:y[99:98];
y[97:97]=(x[97:96]==p)?x[33:32]:y[97:97];
y[95:94]=(x[95:94]==p)?x[31:30]:y[95:94];
y[93:92]=(x[93:92]==p)?x[29:28]:y[93:92];
y[91:90]=(x[91:90]==p)?x[27:26]:y[91:90];
y[89:88]=(x[89:88]==p)?x[25:24]:y[89:88];
y[87:86]=(x[87:86]==p)?x[23:22]:y[87:86];
y[85:84]=(x[85:84]==p)?x[21:20]:y[85:84];
y[83:82]=(x[83:82]==p)?x[19:18]:y[83:82];
y[81:80]=(x[81:80]==p)?x[17:16]:y[81:80];
y[79:78]=(x[79:78]==p)?x[15:14]:y[79:78];
y[77:76]=(x[77:76]==p)?x[13:12]:y[77:76];
y[75:74]=(x[75:74]==p)?x[11:10]:y[75:74];
y[73:72]=(x[73:72]==p)?x[9:8]:y[73:72];
y[71:70]=(x[71:70]==p)?x[7:6]:y[71:70];
y[69:68]=(x[69:68]==p)?x[5:4]:y[69:68];
y[67:66]=(x[67:66]==p)?x[3:2]:y[67:66];
y[65:64]=(x[65:64]==p)?x[1:0]:y[65:64];
end
endmodule



module findxor(a,b,cin,sum,cout);
input [63:0]a,b;
input [129:0]cin;
output [63:0]sum;
output cout;
wire [129:0]c;
assign c[0]=(cin[1:0]==2'b00)?1'b0:1'b1;
assign c[1]=(cin[3:2]==2'b00)?1'b0:1'b1;
assign c[2]=(cin[5:4]==2'b00)?1'b0:1'b1;
assign c[3]=(cin[7:6]==2'b00)?1'b0:1'b1;
assign c[4]=(cin[9:8]==2'b00)?1'b0:1'b1;
assign c[5]=(cin[11:10]==2'b00)?1'b0:1'b1;
assign c[6]=(cin[13:12]==2'b00)?1'b0:1'b1;
assign c[7]=(cin[15:14]==2'b00)?1'b0:1'b1;
assign c[8]=(cin[17:16]==2'b00)?1'b0:1'b1;
assign c[9]=(cin[19:18]==2'b00)?1'b0:1'b1;
assign c[10]=(cin[21:20]==2'b00)?1'b0:1'b1;
assign c[11]=(cin[23:22]==2'b00)?1'b0:1'b1;
assign c[12]=(cin[25:24]==2'b00)?1'b0:1'b1;
assign c[13]=(cin[27:26]==2'b00)?1'b0:1'b1;
assign c[14]=(cin[29:28]==2'b00)?1'b0:1'b1;
assign c[15]=(cin[31:30]==2'b00)?1'b0:1'b1;
assign c[16]=(cin[33:32]==2'b00)?1'b0:1'b1;
assign c[17]=(cin[35:34]==2'b00)?1'b0:1'b1;
assign c[18]=(cin[37:36]==2'b00)?1'b0:1'b1;
assign c[19]=(cin[39:38]==2'b00)?1'b0:1'b1;
assign c[20]=(cin[41:40]==2'b00)?1'b0:1'b1;
assign c[21]=(cin[43:42]==2'b00)?1'b0:1'b1;
assign c[22]=(cin[45:44]==2'b00)?1'b0:1'b1;
assign c[23]=(cin[47:46]==2'b00)?1'b0:1'b1;
assign c[24]=(cin[49:48]==2'b00)?1'b0:1'b1;
assign c[25]=(cin[51:50]==2'b00)?1'b0:1'b1;
assign c[26]=(cin[53:52]==2'b00)?1'b0:1'b1;
assign c[27]=(cin[55:54]==2'b00)?1'b0:1'b1;
assign c[28]=(cin[57:56]==2'b00)?1'b0:1'b1;
assign c[29]=(cin[59:58]==2'b00)?1'b0:1'b1;
assign c[30]=(cin[61:60]==2'b00)?1'b0:1'b1;
assign c[31]=(cin[63:62]==2'b00)?1'b0:1'b1;
assign c[32]=(cin[65:64]==2'b00)?1'b0:1'b1;
assign c[33]=(cin[67:66]==2'b00)?1'b0:1'b1;
assign c[34]=(cin[69:68]==2'b00)?1'b0:1'b1;
assign c[35]=(cin[71:70]==2'b00)?1'b0:1'b1;
assign c[36]=(cin[73:72]==2'b00)?1'b0:1'b1;
assign c[37]=(cin[75:74]==2'b00)?1'b0:1'b1;
assign c[38]=(cin[77:76]==2'b00)?1'b0:1'b1;
assign c[39]=(cin[79:78]==2'b00)?1'b0:1'b1;
assign c[40]=(cin[81:80]==2'b00)?1'b0:1'b1;
assign c[41]=(cin[83:82]==2'b00)?1'b0:1'b1;
assign c[42]=(cin[85:84]==2'b00)?1'b0:1'b1;
assign c[43]=(cin[87:86]==2'b00)?1'b0:1'b1;
assign c[44]=(cin[89:88]==2'b00)?1'b0:1'b1;
assign c[45]=(cin[91:90]==2'b00)?1'b0:1'b1;
assign c[46]=(cin[93:92]==2'b00)?1'b0:1'b1;
assign c[47]=(cin[95:94]==2'b00)?1'b0:1'b1;
assign c[48]=(cin[97:96]==2'b00)?1'b0:1'b1;
assign c[49]=(cin[99:98]==2'b00)?1'b0:1'b1;
assign c[50]=(cin[101:100]==2'b00)?1'b0:1'b1;
assign c[51]=(cin[103:102]==2'b00)?1'b0:1'b1;
assign c[52]=(cin[105:104]==2'b00)?1'b0:1'b1;
assign c[53]=(cin[107:106]==2'b00)?1'b0:1'b1;
assign c[54]=(cin[109:108]==2'b00)?1'b0:1'b1;
assign c[55]=(cin[111:110]==2'b00)?1'b0:1'b1;
assign c[56]=(cin[113:112]==2'b00)?1'b0:1'b1;
assign c[57]=(cin[115:114]==2'b00)?1'b0:1'b1;
assign c[58]=(cin[117:116]==2'b00)?1'b0:1'b1;
assign c[59]=(cin[119:118]==2'b00)?1'b0:1'b1;
assign c[60]=(cin[121:120]==2'b00)?1'b0:1'b1;
assign c[61]=(cin[123:122]==2'b00)?1'b0:1'b1;
assign c[62]=(cin[125:124]==2'b00)?1'b0:1'b1;
assign c[63]=(cin[127:126]==2'b00)?1'b0:1'b1;

xor xor0(sum[0],a[0],b[0],c[0]);
xor xor1(sum[1],a[1],b[1],c[1]);
xor xor2(sum[2],a[2],b[2],c[2]);
xor xor3(sum[3],a[3],b[3],c[3]);
xor xor4(sum[4],a[4],b[4],c[4]);
xor xor5(sum[5],a[5],b[5],c[5]);
xor xor6(sum[6],a[6],b[6],c[6]);
xor xor7(sum[7],a[7],b[7],c[7]);
xor xor8(sum[8],a[8],b[8],c[8]);
xor xor9(sum[9],a[9],b[9],c[9]);
xor xor10(sum[10],a[10],b[10],c[10]);
xor xor11(sum[11],a[11],b[11],c[11]);
xor xor12(sum[12],a[12],b[12],c[12]);
xor xor13(sum[13],a[13],b[13],c[13]);
xor xor14(sum[14],a[14],b[14],c[14]);
xor xor15(sum[15],a[15],b[15],c[15]);
xor xor16(sum[16],a[16],b[16],c[16]);
xor xor17(sum[17],a[17],b[17],c[17]);
xor xor18(sum[18],a[18],b[18],c[18]);
xor xor19(sum[19],a[19],b[19],c[19]);
xor xor20(sum[20],a[20],b[20],c[20]);
xor xor21(sum[21],a[21],b[21],c[21]);
xor xor22(sum[22],a[22],b[22],c[22]);
xor xor23(sum[23],a[23],b[23],c[23]);
xor xor24(sum[24],a[24],b[24],c[24]);
xor xor25(sum[25],a[25],b[25],c[25]);
xor xor26(sum[26],a[26],b[26],c[26]);
xor xor27(sum[27],a[27],b[27],c[27]);
xor xor28(sum[28],a[28],b[28],c[28]);
xor xor29(sum[29],a[29],b[29],c[29]);
xor xor30(sum[30],a[30],b[30],c[30]);
xor xor31(sum[31],a[31],b[31],c[31]);
xor xor32(sum[32],a[32],b[32],c[32]);
xor xor33(sum[33],a[33],b[33],c[33]);
xor xor34(sum[34],a[34],b[34],c[34]);
xor xor35(sum[35],a[35],b[35],c[35]);
xor xor36(sum[36],a[36],b[36],c[36]);
xor xor37(sum[37],a[37],b[37],c[37]);
xor xor38(sum[38],a[38],b[38],c[38]);
xor xor39(sum[39],a[39],b[39],c[39]);
xor xor40(sum[40],a[40],b[40],c[40]);
xor xor41(sum[41],a[41],b[41],c[41]);
xor xor42(sum[42],a[42],b[42],c[42]);
xor xor43(sum[43],a[43],b[43],c[43]);
xor xor44(sum[44],a[44],b[44],c[44]);
xor xor45(sum[45],a[45],b[45],c[45]);
xor xor46(sum[46],a[46],b[46],c[46]);
xor xor47(sum[47],a[47],b[47],c[47]);
xor xor48(sum[48],a[48],b[48],c[48]);
xor xor49(sum[49],a[49],b[49],c[49]);
xor xor50(sum[50],a[50],b[50],c[50]);
xor xor51(sum[51],a[51],b[51],c[51]);
xor xor52(sum[52],a[52],b[52],c[52]);
xor xor53(sum[53],a[53],b[53],c[53]);
xor xor54(sum[54],a[54],b[54],c[54]);
xor xor55(sum[55],a[55],b[55],c[55]);
xor xor56(sum[56],a[56],b[56],c[56]);
xor xor57(sum[57],a[57],b[57],c[57]);
xor xor58(sum[58],a[58],b[58],c[58]);
xor xor59(sum[59],a[59],b[59],c[59]);
xor xor60(sum[60],a[60],b[60],c[60]);
xor xor61(sum[61],a[61],b[61],c[61]);
xor xor62(sum[62],a[62],b[62],c[62]);
xor xor63(sum[63],a[63],b[63],c[63]);
assign cout=c[64];
endmodule

